package shared_pkg;
    int error_count = 0;
    int correct_count = 0;

    logic test_finished;
endpackage